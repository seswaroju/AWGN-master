`timescale 1ns / 1ps
//------------------------------------------------------------------------------
//
// cos_table.v
//
// This file is part of the AWGN IP core
//
// Description
//     Coefficients ROM table for cosine polynomial degree 1.
//
//------------------------------------------------------------------------------


module cos_table(
    // System signals
    input clock,
    
    // Data interface
    input [6:0] addr,       //read address
    output reg [11:0] c1,   // coefficient c1
    output reg [18:0] c0    // coefficient c0
    );
    
    // local variables
    reg [30:0] d;       // {c1, c0}
    
    //Table 
    always @(*) begin
        case (addr)
		7'd0 : d = 31'b000000011001_10000000000000000110;
		7'd1 : d = 31'b000001001011_10000000000001010101;
		7'd2 : d = 31'b000001111101_10000000000011110011;
		7'd3 : d = 31'b000010101111_10000000000111100000;
		7'd4 : d = 31'b000011100010_10000000001100011011;
		7'd5 : d = 31'b000100010100_10000000010010100101;
		7'd6 : d = 31'b000101000110_10000000011001111101;
		7'd7 : d = 31'b000101111000_10000000100010100100;
		7'd8 : d = 31'b000110101010_10000000101100011001;
		7'd9 : d = 31'b000111011100_10000000110111011011;
		7'd10 : d = 31'b001000001110_10000001000011101011;
		7'd11 : d = 31'b001001000000_10000001010001000111;
		7'd12 : d = 31'b001001110001_10000001011111110000;
		7'd13 : d = 31'b001010100011_10000001101111100110;
		7'd14 : d = 31'b001011010101_10000010000000100111;
		7'd15 : d = 31'b001100000110_10000010010010110011;
		7'd16 : d = 31'b001100110111_10000010100110001010;
		7'd17 : d = 31'b001101101000_10000010111010101011;
		7'd18 : d = 31'b001110011001_10000011010000010110;
		7'd19 : d = 31'b001111001010_10000011100111001010;
		7'd20 : d = 31'b001111111011_10000011111111000101;
		7'd21 : d = 31'b010000101100_10000100011000001001;
		7'd22 : d = 31'b010001011100_10000100110010010011;
		7'd23 : d = 31'b010010001100_10000101001101100011;
		7'd24 : d = 31'b010010111101_10000101101001111000;
		7'd25 : d = 31'b010011101100_10000110000111010010;
		7'd26 : d = 31'b010100011100_10000110100101101111;
		7'd27 : d = 31'b010101001100_10000111000101001111;
		7'd28 : d = 31'b010101111011_10000111100101110000;
		7'd29 : d = 31'b010110101010_10001000000111010011;
		7'd30 : d = 31'b010111011001_10001000101001110101;
		7'd31 : d = 31'b011000001000_10001001001101010101;
		7'd32 : d = 31'b011000110110_10001001110001110100;
		7'd33 : d = 31'b011001100100_10001010010111001110;
		7'd34 : d = 31'b011010010010_10001010111101100100;
		7'd35 : d = 31'b011011000000_10001011100100110101;
		7'd36 : d = 31'b011011101101_10001100001100111110;
		7'd37 : d = 31'b011100011011_10001100110110000000;
		7'd38 : d = 31'b011101001000_10001101011111111000;
		7'd39 : d = 31'b011101110100_10001110001010100101;
		7'd40 : d = 31'b011110100000_10001110110110000110;
		7'd41 : d = 31'b011111001100_10001111100010011010;
		7'd42 : d = 31'b011111111000_10010000001111011111;
		7'd43 : d = 31'b0100000100100_10010000111101010101;
		7'd44 : d = 31'b0100001001111_10010001101011111001;
		7'd45 : d = 31'b0100001111010_10010010011011001001;
		7'd46 : d = 31'b0100010100100_10010011001011000110;
		7'd47 : d = 31'b0100011001110_10010011111011101100;
		7'd48 : d = 31'b0100011111000_10010100101100111100;
		7'd49 : d = 31'b0100100100001_10010101011110110010;
		7'd50 : d = 31'b0100101001011_10010110010001001101;
		7'd51 : d = 31'b0100101110011_10010111000100001101;
		7'd52 : d = 31'b0100110011100_10010111110111101110;
		7'd53 : d = 31'b0100111000100_10011000101011110001;
		7'd54 : d = 31'b0100111101011_10011001100000010010;
		7'd55 : d = 31'b0101000010010_10011010010101010000;
		7'd56 : d = 31'b0101000111001_10011011001010101010;
		7'd57 : d = 31'b0101001100000_10011100000000011110;
		7'd58 : d = 31'b0101010000110_10011100110110101001;
		7'd59 : d = 31'b0101010101100_10011101101101001011;
		7'd60 : d = 31'b0101011010001_10011110100100000001;
		7'd61 : d = 31'b0101011110110_10011111011011001010;
		7'd62 : d = 31'b0101100011010_10100000010010100011;
		7'd63 : d = 31'b0101100111110_10100001001010001011;
		7'd64 : d = 31'b0101101100010_10100010000010000000;
		7'd65 : d = 31'b0101110000101_10100010111010000001;
		7'd66 : d = 31'b0101110100111_10100011110010001010;
		7'd67 : d = 31'b0101111001001_10100100101010011010;
		7'd68 : d = 31'b0101111101011_10100101100010110000;
		7'd69 : d = 31'b0110000001101_10100110011011001000;
		7'd70 : d = 31'b0110000101101_10100111010011100010;
		7'd71 : d = 31'b0110001001110_10101000001011111100;
		7'd72 : d = 31'b0110001101110_10101001000100010010;
		7'd73 : d = 31'b0110010001101_10101001111100100100;
		7'd74 : d = 31'b0110010101100_10101010110100101110;
		7'd75 : d = 31'b0110011001010_10101011101100110000;
		7'd76 : d = 31'b0110011101000_10101100100100100110;
		7'd77 : d = 31'b0110100000110_10101101011100010000;
		7'd78 : d = 31'b0110100100011_10101110010011101010;
		7'd79 : d = 31'b0110100111111_10101111001010110010;
		7'd80 : d = 31'b0110101011011_10110000000001101000;
		7'd81 : d = 31'b0110101110110_10110000111000000111;
		7'd82 : d = 31'b0110110010001_10110001101110001111;
		7'd83 : d = 31'b0110110101100_10110010100011111101;
		7'd84 : d = 31'b0110111000110_10110011011001001110;
		7'd85 : d = 31'b0110111011111_10110100001110000010;
		7'd86 : d = 31'b0110111111000_10110101000010010100;
		7'd87 : d = 31'b0111000010000_10110101110110000101;
		7'd88 : d = 31'b0111000101000_10110110101001010000;
		7'd89 : d = 31'b0111000111111_10110111011011110100;
		7'd90 : d = 31'b0111001010101_10111000001101101111;
		7'd91 : d = 31'b0111001101011_10111000111110111110;
		7'd92 : d = 31'b0111010000001_10111001101111100000;
		7'd93 : d = 31'b0111010010110_10111010011111010010;
		7'd94 : d = 31'b0111010101010_10111011001110010001;
		7'd95 : d = 31'b0111010111110_10111011111100011101;
		7'd96 : d = 31'b0111011010001_10111100101001110001;
		7'd97 : d = 31'b0111011100100_10111101010110001101;
		7'd98 : d = 31'b0111011110110_10111110000001101110;
		7'd99 : d = 31'b0111100001000_10111110101100010001;
		7'd100 : d = 31'b0111100011000_10111111010101110101;
		7'd101 : d = 31'b0111100101001_10111111111110010111;
		7'd102 : d = 31'b0111100111001_11000000100101110101;
		7'd103 : d = 31'b0111101001000_11000001001100001101;
		7'd104 : d = 31'b0111101010110_11000001110001011101;
		7'd105 : d = 31'b0111101100100_11000010010101100010;
		7'd106 : d = 31'b0111101110010_11000010111000011010;
		7'd107 : d = 31'b0111101111111_11000011011010000011;
		7'd108 : d = 31'b0111110001011_11000011111010011011;
		7'd109 : d = 31'b0111110010110_11000100011001011111;
		7'd110 : d = 31'b0111110100001_11000100110111001110;
		7'd111 : d = 31'b0111110101100_11000101010011100101;
		7'd112 : d = 31'b0111110110110_11000101101110100011;
		7'd113 : d = 31'b0111110111111_11000110001000000100;
		7'd114 : d = 31'b0111111000111_11000110100000000110;
		7'd115 : d = 31'b0111111001111_11000110110110101001;
		7'd116 : d = 31'b0111111010111_11000111001011101001;
		7'd117 : d = 31'b0111111011110_11000111011111000100;
		7'd118 : d = 31'b0111111100100_11000111110000111000;
		7'd119 : d = 31'b0111111101001_11001000000001000100;
		7'd120 : d = 31'b0111111101110_11001000001111100100;
		7'd121 : d = 31'b0111111110010_11001000011100011000;
		7'd122 : d = 31'b0111111110110_11001000100111011100;
		7'd123 : d = 31'b0111111111001_11001000110000110000;
		7'd124 : d = 31'b0111111111100_11001000111000010000;
		7'd125 : d = 31'b0111111111110_11001000111101111011;
		7'd126 : d = 31'b0111111111111_11001001000001110000;
		7'd127 : d = 31'b0111111111111_11001001000011101011;
        	default: d = 31'd0;
        endcase
    end
    
    // Output Data
    always @(posedge clock) begin
        c1 <= d[30:19];
        c0 <= d[18:0];
    end    
endmodule
