`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//
//	log_coeff_table.v
//
//	Description: This module is used as a rom for generating coeffs for log function.
// 
//////////////////////////////////////////////////////////////////////////////////


module log_coeff_table(
    input clock,
    // Data Interface
    input [7:0] log_addr,
    output reg [12:0] log_c2,
    output reg [21:0] log_c1,
    output reg [29:0] log_c0
    );
    
    // Local Variables
    reg [64:0] d;
    
    //Table
    always @(*) begin
        case (log_addr)
			8'd0 : d = 65'b1001101110101_1011110011001100001000_100000000011110011001100001000;
        8'd1 : d = 65'b1001101001110_1011110001010011000000_100000000011110001010011000000;
        8'd2 : d = 65'b1001100101000_1011101111011010110100_100000000011101111011010110100;
        8'd3 : d = 65'b1001100000010_1011101101100011100011_100000000011101101100011100011;
        8'd4 : d = 65'b1001011011101_1011101011101101001101_100000000011101011101101001101;
        8'd5 : d = 65'b1001010111000_1011101001110111110001_100000000011101001110111110001;
        8'd6 : d = 65'b1001010010011_1011101000000011001110_100000000011101000000011001110;
        8'd7 : d = 65'b1001001101111_1011100110001111100100_100000000011100110001111100100;
        8'd8 : d = 65'b1001001001100_1011100100011100110010_100000000011100100011100110010;
        8'd9 : d = 65'b1001000101001_1011100010101010110111_100000000011100010101010110111;
        8'd10 : d = 65'b1001000000110_1011100000111001110011_100000000011100000111001110011;
        8'd11 : d = 65'b1000111100011_1011011111001001100101_100000000011011111001001100101;
        8'd12 : d = 65'b1000111000001_1011011101011010001100_100000000011011101011010001100;
        8'd13 : d = 65'b1000110100000_1011011011101011101001_100000000011011011101011101001;
        8'd14 : d = 65'b1000101111110_1011011001111101111001_100000000011011001111101111001;
        8'd15 : d = 65'b1000101011101_1011011000010000111110_100000000011011000010000111110;
        8'd16 : d = 65'b1000100111101_1011010110100100110101_100000000011010110100100110101;
        8'd17 : d = 65'b1000100011101_1011010100111001011111_100000000011010100111001011111;
        8'd18 : d = 65'b1000011111101_1011010011001110111011_100000000011010011001110111011;
        8'd19 : d = 65'b1000011011101_1011010001100101001001_100000000011010001100101001001;
        8'd20 : d = 65'b1000010111110_1011001111111100001000_100000000011001111111100001000;
        8'd21 : d = 65'b1000010011111_1011001110010011110111_100000000011001110010011110111;
        8'd22 : d = 65'b1000010000001_1011001100101100010110_100000000011001100101100010110;
        8'd23 : d = 65'b1000001100011_1011001011000101100100_100000000011001011000101100100;
        8'd24 : d = 65'b1000001000101_1011001001011111100010_100000000011001001011111100010;
        8'd25 : d = 65'b1000000100111_1011000111111010001110_100000000011000111111010001110;
        8'd26 : d = 65'b1000000001010_1011000110010101100111_100000000011000110010101100111;
        8'd27 : d = 65'b0111111101101_1011000100110001101110_100000000011000100110001101110;
        8'd28 : d = 65'b0111111010000_1011000011001110100010_100000000011000011001110100010;
        8'd29 : d = 65'b0111110110100_1011000001101100000011_100000000011000001101100000011;
        8'd30 : d = 65'b0111110011000_1011000000001010001111_100000000011000000001010001111;
        8'd31 : d = 65'b0111101111100_1010111110101001000111_100000000010111110101001000111;
        8'd32 : d = 65'b0111101100001_1010111101001000101010_100000000010111101001000101010;
        8'd33 : d = 65'b0111101000110_1010111011101000111000_100000000010111011101000111000;
        8'd34 : d = 65'b0111100101011_1010111010001001110000_100000000010111010001001110000;
        8'd35 : d = 65'b0111100010000_1010111000101011010010_100000000010111000101011010010;
        8'd36 : d = 65'b0111011110110_1010110111001101011101_100000000010110111001101011101;
        8'd37 : d = 65'b0111011011100_1010110101110000010001_100000000010110101110000010001;
        8'd38 : d = 65'b0111011000010_1010110100010011101110_100000000010110100010011101110;
        8'd39 : d = 65'b0111010101001_1010110010110111110010_100000000010110010110111110010;
        8'd40 : d = 65'b0111010001111_1010110001011100011110_100000000010110001011100011110;
        8'd41 : d = 65'b0111001110110_1010110000000001110010_100000000010110000000001110010;
        8'd42 : d = 65'b0111001011110_1010101110100111101100_100000000010101110100111101100;
        8'd43 : d = 65'b0111001000101_1010101101001110001101_100000000010101101001110001101;
        8'd44 : d = 65'b0111000101101_1010101011110101010100_100000000010101011110101010100;
        8'd45 : d = 65'b0111000010101_1010101010011101000001_100000000010101010011101000001;
        8'd46 : d = 65'b0110111111101_1010101001000101010011_100000000010101001000101010011;
        8'd47 : d = 65'b0110111100101_1010100111101110001011_100000000010100111101110001011;
        8'd48 : d = 65'b0110111001110_1010100110010111100110_100000000010100110010111100110;
        8'd49 : d = 65'b0110110110111_1010100101000001100111_100000000010100101000001100111;
        8'd50 : d = 65'b0110110100000_1010100011101100001011_100000000010100011101100001011;
        8'd51 : d = 65'b0110110001001_1010100010010111010010_100000000010100010010111010010;
        8'd52 : d = 65'b0110101110011_1010100001000010111101_100000000010100001000010111101;
        8'd53 : d = 65'b0110101011101_1010011111101111001010_100000000010011111101111001010;
        8'd54 : d = 65'b0110101000111_1010011110011011111011_100000000010011110011011111011;
        8'd55 : d = 65'b0110100110001_1010011101001001001101_100000000010011101001001001101;
        8'd56 : d = 65'b0110100011011_1010011011110111000001_100000000010011011110111000001;
        8'd57 : d = 65'b0110100000110_1010011010100101010111_100000000010011010100101010111;
        8'd58 : d = 65'b0110011110001_1010011001010100001110_100000000010011001010100001110;
        8'd59 : d = 65'b0110011011100_1010011000000011100110_100000000010011000000011100110;
        8'd60 : d = 65'b0110011000111_1010010110110011011111_100000000010010110110011011111;
        8'd61 : d = 65'b0110010110011_1010010101100011111000_100000000010010101100011111000;
        8'd62 : d = 65'b0110010011110_1010010100010100110001_100000000010010100010100110001;
        8'd63 : d = 65'b0110010001010_1010010011000110001001_100000000010010011000110001001;
        8'd64 : d = 65'b0110001110110_1010010001111000000001_100000000010010001111000000001;
        8'd65 : d = 65'b0110001100010_1010010000101010011000_100000000010010000101010011000;
        8'd66 : d = 65'b0110001001111_1010001111011101001110_100000000010001111011101001110;
        8'd67 : d = 65'b0110000111011_1010001110010000100011_100000000010001110010000100011;
        8'd68 : d = 65'b0110000101000_1010001101000100010101_100000000010001101000100010101;
        8'd69 : d = 65'b0110000010101_1010001011111000100110_100000000010001011111000100110;
        8'd70 : d = 65'b0110000000010_1010001010101101010100_100000000010001010101101010100;
        8'd71 : d = 65'b0101111101111_1010001001100010100000_100000000010001001100010100000;
        8'd72 : d = 65'b0101111011101_1010001000011000001001_100000000010001000011000001001;
        8'd73 : d = 65'b0101111001010_1010000111001110001111_100000000010000111001110001111;
        8'd74 : d = 65'b0101110111000_1010000110000100110001_100000000010000110000100110001;
        8'd75 : d = 65'b0101110100110_1010000100111011110000_100000000010000100111011110000;
        8'd76 : d = 65'b0101110010100_1010000011110011001011_100000000010000011110011001011;
        8'd77 : d = 65'b0101110000010_1010000010101011000001_100000000010000010101011000001;
        8'd78 : d = 65'b0101101110001_1010000001100011010100_100000000010000001100011010100;
        8'd79 : d = 65'b0101101011111_1010000000011100000010_100000000010000000011100000010;
        8'd80 : d = 65'b0101101001110_1001111111010101001010_100000000001111111010101001010;
        8'd81 : d = 65'b0101100111101_1001111110001110101110_100000000001111110001110101110;
        8'd82 : d = 65'b0101100101100_1001111101001000101100_100000000001111101001000101100;
        8'd83 : d = 65'b0101100011011_1001111100000011000101_100000000001111100000011000101;
        8'd84 : d = 65'b0101100001010_1001111010111101111000_100000000001111010111101111000;
        8'd85 : d = 65'b0101011111010_1001111001111001000101_100000000001111001111001000101;
        8'd86 : d = 65'b0101011101001_1001111000110100101100_100000000001111000110100101100;
        8'd87 : d = 65'b0101011011001_1001110111110000101100_100000000001110111110000101100;
        8'd88 : d = 65'b0101011001001_1001110110101101000101_100000000001110110101101000101;
        8'd89 : d = 65'b0101010111001_1001110101101001110111_100000000001110101101001110111;
        8'd90 : d = 65'b0101010101001_1001110100100111000010_100000000001110100100111000010;
        8'd91 : d = 65'b0101010011010_1001110011100100100110_100000000001110011100100100110;
        8'd92 : d = 65'b0101010001010_1001110010100010100010_100000000001110010100010100010;
        8'd93 : d = 65'b0101001111011_1001110001100000110111_100000000001110001100000110111;
        8'd94 : d = 65'b0101001101011_1001110000011111100011_100000000001110000011111100011;
        8'd95 : d = 65'b0101001011100_1001101111011110100111_100000000001101111011110100111;
        8'd96 : d = 65'b0101001001101_1001101110011110000011_100000000001101110011110000011;
        8'd97 : d = 65'b0101000111110_1001101101011101110110_100000000001101101011101110110;
        8'd98 : d = 65'b0101000101111_1001101100011110000001_100000000001101100011110000001;
        8'd99 : d = 65'b0101000100001_1001101011011110100010_100000000001101011011110100010;
        8'd100 : d = 65'b0101000010010_1001101010011111011010_100000000001101010011111011010;
        8'd101 : d = 65'b0101000000100_1001101001100000101001_100000000001101001100000101001;
        8'd102 : d = 65'b0100111110110_1001101000100010001110_100000000001101000100010001110;
        8'd103 : d = 65'b0100111100111_1001100111100100001001_100000000001100111100100001001;
        8'd104 : d = 65'b0100111011001_1001100110100110011011_100000000001100110100110011011;
        8'd105 : d = 65'b0100111001011_1001100101101001000010_100000000001100101101001000010;
        8'd106 : d = 65'b0100110111110_1001100100101011111111_100000000001100100101011111111;
        8'd107 : d = 65'b0100110110000_1001100011101111010001_100000000001100011101111010001;
        8'd108 : d = 65'b0100110100010_1001100010110010111001_100000000001100010110010111001;
        8'd109 : d = 65'b0100110010101_1001100001110110110110_100000000001100001110110110110;
        8'd110 : d = 65'b0100110001000_1001100000111011000111_100000000001100000111011000111;
        8'd111 : d = 65'b0100101111010_1001011111111111101110_100000000001011111111111101110;
        8'd112 : d = 65'b0100101101101_1001011111000100101001_100000000001011111000100101001;
        8'd113 : d = 65'b0100101100000_1001011110001001111001_100000000001011110001001111001;
        8'd114 : d = 65'b0100101010011_1001011101001111011101_100000000001011101001111011101;
        8'd115 : d = 65'b0100101000110_1001011100010101010101_100000000001011100010101010101;
        8'd116 : d = 65'b0100100111010_1001011011011011100001_100000000001011011011011100001;
        8'd117 : d = 65'b0100100101101_1001011010100010000001_100000000001011010100010000001;
        8'd118 : d = 65'b0100100100000_1001011001101000110101_100000000001011001101000110101;
        8'd119 : d = 65'b0100100010100_1001011000101111111100_100000000001011000101111111100;
        8'd120 : d = 65'b0100100001000_1001010111110111010111_100000000001010111110111010111;
        8'd121 : d = 65'b0100011111011_1001010110111111000100_100000000001010110111111000100;
        8'd122 : d = 65'b0100011101111_1001010110000111000101_100000000001010110000111000101;
        8'd123 : d = 65'b0100011100011_1001010101001111011000_100000000001010101001111011000;
        8'd124 : d = 65'b0100011010111_1001010100010111111111_100000000001010100010111111111;
        8'd125 : d = 65'b0100011001011_1001010011100000111000_100000000001010011100000111000;
        8'd126 : d = 65'b0100011000000_1001010010101010000011_100000000001010010101010000011;
        8'd127 : d = 65'b0100010110100_1001010001110011100000_100000000001010001110011100000;
        8'd128 : d = 65'b0100010101000_1001010000111101010000_100000000001010000111101010000;
        8'd129 : d = 65'b0100010011101_1001010000000111010010_100000000001010000000111010010;
        8'd130 : d = 65'b0100010010010_1001001111010001100110_100000000001001111010001100110;
        8'd131 : d = 65'b0100010000110_1001001110011100001011_100000000001001110011100001011;
        8'd132 : d = 65'b0100001111011_1001001101100111000010_100000000001001101100111000010;
        8'd133 : d = 65'b0100001110000_1001001100110010001010_100000000001001100110010001010;
        8'd134 : d = 65'b0100001100101_1001001011111101100100_100000000001001011111101100100;
        8'd135 : d = 65'b0100001011010_1001001011001001001111_100000000001001011001001001111;
        8'd136 : d = 65'b0100001001111_1001001010010101001011_100000000001001010010101001011;
        8'd137 : d = 65'b0100001000100_1001001001100001011000_100000000001001001100001011000;
        8'd138 : d = 65'b0100000111010_1001001000101101110110_100000000001001000101101110110;
        8'd139 : d = 65'b0100000101111_1001000111111010100101_100000000001000111111010100101;
        8'd140 : d = 65'b0100000100100_1001000111000111100100_100000000001000111000111100100;
        8'd141 : d = 65'b0100000011010_1001000110010100110011_100000000001000110010100110011;
        8'd142 : d = 65'b0100000001111_1001000101100010010011_100000000001000101100010010011;
        8'd143 : d = 65'b0100000000101_1001000100110000000011_100000000001000100110000000011;
        8'd144 : d = 65'b0011111111011_1001000011111110000011_100000000001000011111110000011;
        8'd145 : d = 65'b0011111110001_1001000011001100010011_100000000001000011001100010011;
        8'd146 : d = 65'b0011111100111_1001000010011010110010_100000000001000010011010110010;
        8'd147 : d = 65'b0011111011101_1001000001101001100010_100000000001000001101001100010;
        8'd148 : d = 65'b0011111010011_1001000000111000100001_100000000001000000111000100001;
        8'd149 : d = 65'b0011111001001_1001000000000111101111_100000000001000000000111101111;
        8'd150 : d = 65'b0011110111111_1000111111010111001101_100000000000111111010111001101;
        8'd151 : d = 65'b0011110110101_1000111110100110111010_100000000000111110100110111010;
        8'd152 : d = 65'b0011110101100_1000111101110110110111_100000000000111101110110110111;
        8'd153 : d = 65'b0011110100010_1000111101000111000010_100000000000111101000111000010;
        8'd154 : d = 65'b0011110011001_1000111100010111011100_100000000000111100010111011100;
        8'd155 : d = 65'b0011110001111_1000111011101000000101_100000000000111011101000000101;
        8'd156 : d = 65'b0011110000110_1000111010111000111101_100000000000111010111000111101;
        8'd157 : d = 65'b0011101111100_1000111010001010000011_100000000000111010001010000011;
        8'd158 : d = 65'b0011101110011_1000111001011011011000_100000000000111001011011011000;
        8'd159 : d = 65'b0011101101010_1000111000101100111011_100000000000111000101100111011;
        8'd160 : d = 65'b0011101100001_1000110111111110101100_100000000000110111111110101100;
        8'd161 : d = 65'b0011101011000_1000110111010000101100_100000000000110111010000101100;
        8'd162 : d = 65'b0011101001111_1000110110100010111010_100000000000110110100010111010;
        8'd163 : d = 65'b0011101000110_1000110101110101010101_100000000000110101110101010101;
        8'd164 : d = 65'b0011100111101_1000110101000111111111_100000000000110101000111111111;
        8'd165 : d = 65'b0011100110100_1000110100011010110110_100000000000110100011010110110;
        8'd166 : d = 65'b0011100101100_1000110011101101111011_100000000000110011101101111011;
        8'd167 : d = 65'b0011100100011_1000110011000001001101_100000000000110011000001001101;
        8'd168 : d = 65'b0011100011010_1000110010010100101101_100000000000110010010100101101;
        8'd169 : d = 65'b0011100010010_1000110001101000011011_100000000000110001101000011011;
        8'd170 : d = 65'b0011100001001_1000110000111100010101_100000000000110000111100010101;
        8'd171 : d = 65'b0011100000001_1000110000010000011101_100000000000110000010000011101;
        8'd172 : d = 65'b0011011111001_1000101111100100110010_100000000000101111100100110010;
        8'd173 : d = 65'b0011011110000_1000101110111001010100_100000000000101110111001010100;
        8'd174 : d = 65'b0011011101000_1000101110001110000011_100000000000101110001110000011;
        8'd175 : d = 65'b0011011100000_1000101101100010111111_100000000000101101100010111111;
        8'd176 : d = 65'b0011011011000_1000101100111000001000_100000000000101100111000001000;
        8'd177 : d = 65'b0011011010000_1000101100001101011101_100000000000101100001101011101;
        8'd178 : d = 65'b0011011001000_1000101011100010111110_100000000000101011100010111110;
        8'd179 : d = 65'b0011011000000_1000101010111000101101_100000000000101010111000101101;
        8'd180 : d = 65'b0011010111000_1000101010001110100111_100000000000101010001110100111;
        8'd181 : d = 65'b0011010110000_1000101001100100101110_100000000000101001100100101110;
        8'd182 : d = 65'b0011010101000_1000101000111011000001_100000000000101000111011000001;
        8'd183 : d = 65'b0011010100000_1000101000010001100001_100000000000101000010001100001;
        8'd184 : d = 65'b0011010011001_1000100111101000001100_100000000000100111101000001100;
        8'd185 : d = 65'b0011010010001_1000100110111111000011_100000000000100110111111000011;
        8'd186 : d = 65'b0011010001001_1000100110010110000111_100000000000100110010110000111;
        8'd187 : d = 65'b0011010000010_1000100101101101010110_100000000000100101101101010110;
        8'd188 : d = 65'b0011001111010_1000100101000100110000_100000000000100101000100110000;
        8'd189 : d = 65'b0011001110011_1000100100011100010111_100000000000100100011100010111;
        8'd190 : d = 65'b0011001101100_1000100011110100001001_100000000000100011110100001001;
        8'd191 : d = 65'b0011001100100_1000100011001100000111_100000000000100011001100000111;
        8'd192 : d = 65'b0011001011101_1000100010100100010000_100000000000100010100100010000;
        8'd193 : d = 65'b0011001010110_1000100001111100100100_100000000000100001111100100100;
        8'd194 : d = 65'b0011001001111_1000100001010101000011_100000000000100001010101000011;
        8'd195 : d = 65'b0011001000111_1000100000101101101110_100000000000100000101101101110;
        8'd196 : d = 65'b0011001000000_1000100000000110100100_100000000000100000000110100100;
        8'd197 : d = 65'b0011000111001_1000011111011111100101_100000000000011111011111100101;
        8'd198 : d = 65'b0011000110010_1000011110111000110001_100000000000011110111000110001;
        8'd199 : d = 65'b0011000101011_1000011110010010001000_100000000000011110010010001000;
        8'd200 : d = 65'b0011000100100_1000011101101011101010_100000000000011101101011101010;
        8'd201 : d = 65'b0011000011110_1000011101000101010110_100000000000011101000101010110;
        8'd202 : d = 65'b0011000010111_1000011100011111001101_100000000000011100011111001101;
        8'd203 : d = 65'b0011000010000_1000011011111001001111_100000000000011011111001001111;
        8'd204 : d = 65'b0011000001001_1000011011010011011011_100000000000011011010011011011;
        8'd205 : d = 65'b0011000000011_1000011010101101110010_100000000000011010101101110010;
        8'd206 : d = 65'b0010111111100_1000011010001000010011_100000000000011010001000010011;
        8'd207 : d = 65'b0010111110101_1000011001100010111111_100000000000011001100010111111;
        8'd208 : d = 65'b0010111101111_1000011000111101110101_100000000000011000111101110101;
        8'd209 : d = 65'b0010111101000_1000011000011000110101_100000000000011000011000110101;
        8'd210 : d = 65'b0010111100010_1000010111110011111111_100000000000010111110011111111;
        8'd211 : d = 65'b0010111011011_1000010111001111010100_100000000000010111001111010100;
        8'd212 : d = 65'b0010111010101_1000010110101010110010_100000000000010110101010110010;
        8'd213 : d = 65'b0010111001111_1000010110000110011010_100000000000010110000110011010;
        8'd214 : d = 65'b0010111001000_1000010101100010001100_100000000000010101100010001100;
        8'd215 : d = 65'b0010111000010_1000010100111110001000_100000000000010100111110001000;
        8'd216 : d = 65'b0010110111100_1000010100011010001110_100000000000010100011010001110;
        8'd217 : d = 65'b0010110110110_1000010011110110011110_100000000000010011110110011110;
        8'd218 : d = 65'b0010110101111_1000010011010010110111_100000000000010011010010110111;
        8'd219 : d = 65'b0010110101001_1000010010101111011010_100000000000010010101111011010;
        8'd220 : d = 65'b0010110100011_1000010010001100000110_100000000000010010001100000110;
        8'd221 : d = 65'b0010110011101_1000010001101000111100_100000000000010001101000111100;
        8'd222 : d = 65'b0010110010111_1000010001000101111011_100000000000010001000101111011;
        8'd223 : d = 65'b0010110010001_1000010000100011000011_100000000000010000100011000011;
        8'd224 : d = 65'b0010110001011_1000010000000000010101_100000000000010000000000010101;
        8'd225 : d = 65'b0010110000101_1000001111011101110000_100000000000001111011101110000;
        8'd226 : d = 65'b0010110000000_1000001110111011010100_100000000000001110111011010100;
        8'd227 : d = 65'b0010101111010_1000001110011001000010_100000000000001110011001000010;
        8'd228 : d = 65'b0010101110100_1000001101110110111000_100000000000001101110110111000;
        8'd229 : d = 65'b0010101101110_1000001101010100110111_100000000000001101010100110111;
        8'd230 : d = 65'b0010101101000_1000001100110011000000_100000000000001100110011000000;
        8'd231 : d = 65'b0010101100011_1000001100010001010001_100000000000001100010001010001;
        8'd232 : d = 65'b0010101011101_1000001011101111101011_100000000000001011101111101011;
        8'd233 : d = 65'b0010101011000_1000001011001110001110_100000000000001011001110001110;
        8'd234 : d = 65'b0010101010010_1000001010101100111001_100000000000001010101100111001;
        8'd235 : d = 65'b0010101001100_1000001010001011101101_100000000000001010001011101101;
        8'd236 : d = 65'b0010101000111_1000001001101010101010_100000000000001001101010101010;
        8'd237 : d = 65'b0010101000001_1000001001001001110000_100000000000001001001001110000;
        8'd238 : d = 65'b0010100111100_1000001000101000111110_100000000000001000101000111110;
        8'd239 : d = 65'b0010100110111_1000001000001000010100_100000000000001000001000010100;
        8'd240 : d = 65'b0010100110001_1000000111100111110011_100000000000000111100111110011;
        8'd241 : d = 65'b0010100101100_1000000111000111011010_100000000000000111000111011010;
        8'd242 : d = 65'b0010100100111_1000000110100111001010_100000000000000110100111001010;
        8'd243 : d = 65'b0010100100001_1000000110000111000001_100000000000000110000111000001;
        8'd244 : d = 65'b0010100011100_1000000101100111000001_100000000000000101100111000001;
        8'd245 : d = 65'b0010100010111_1000000101000111001010_100000000000000101000111001010;
        8'd246 : d = 65'b0010100010010_1000000100100111011010_100000000000000100100111011010;
        8'd247 : d = 65'b0010100001101_1000000100000111110010_100000000000000100000111110010;
        8'd248 : d = 65'b0010100000111_1000000011101000010011_100000000000000011101000010011;
        8'd249 : d = 65'b0010100000010_1000000011001000111011_100000000000000011001000111011;
        8'd250 : d = 65'b0010011111101_1000000010101001101011_100000000000000010101001101011;
        8'd251 : d = 65'b0010011111000_1000000010001010100011_100000000000000010001010100011;
        8'd252 : d = 65'b0010011110011_1000000001101011100011_100000000000000001101011100011;
        8'd253 : d = 65'b0010011101110_1000000001001100101011_100000000000000001001100101011;
        8'd254 : d = 65'b0010011101001_1000000000101101111011_100000000000000000101101111011;
        8'd255 : d = 65'b0010011100100_1000000000001111010010_100000000000000000001111010010;
        default: d = 65'd0;
        endcase
    end

    // Output Data
    always @(posedge clock) begin
        log_c2 <= d[64:52];
        log_c1 <= d[51:30];
        log_c0 <= d[29:0];
    end  
endmodule
