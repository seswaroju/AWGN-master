`timescale 1ns / 1ps
//------------------------------------------------------------------------------
//
// cos_table.v
//
// This file is part of the AWGN IP core
//
// Description
//     Coefficients ROM table for cosine polynomial degree 1.
//
//------------------------------------------------------------------------------


module cos_table(
    // System signals
    input clock,
    
    // Data interface
    input [6:0] addr,       //read address
    output reg [11:0] c1,   // coefficient c1
    output reg [18:0] c0    // coefficient c0
    );
    
    // local variables
    reg [30:0] d;       // {c1, c0}
    
    //Table 
    always @(*) begin
        case (addr)
		7'd0 : d = 31'b000000000110_1000000000000000001;
        7'd1 : d = 31'b000000010010_1000000000000010000;
        7'd2 : d = 31'b000000011111_1000000000000101110;
        7'd3 : d = 31'b000000101011_1000000000001011100;
        7'd4 : d = 31'b000000110111_1000000000010011000;
        7'd5 : d = 31'b000001000011_1000000000011100011;
        7'd6 : d = 31'b000001010000_1000000000100111101;
        7'd7 : d = 31'b000001011100_1000000000110100110;
        7'd8 : d = 31'b000001101000_1000000001000011110;
        7'd9 : d = 31'b000001110100_1000000001010100101;
        7'd10 : d = 31'b000010000000_1000000001100111010;
        7'd11 : d = 31'b000010001101_1000000001111011110;
        7'd12 : d = 31'b000010011001_1000000010010010001;
        7'd13 : d = 31'b000010100101_1000000010101010010;
        7'd14 : d = 31'b000010110001_1000000011000100010;
        7'd15 : d = 31'b000010111101_1000000011100000000;
        7'd16 : d = 31'b000011001001_1000000011111101100;
        7'd17 : d = 31'b000011010101_1000000100011100111;
        7'd18 : d = 31'b000011100001_1000000100111101111;
        7'd19 : d = 31'b000011101101_1000000101100000110;
        7'd20 : d = 31'b000011111001_1000000110000101010;
        7'd21 : d = 31'b000100000101_1000000110101011100;
        7'd22 : d = 31'b000100010001_1000000111010011011;
        7'd23 : d = 31'b000100011100_1000000111111101000;
        7'd24 : d = 31'b000100101000_1000001000101000010;
        7'd25 : d = 31'b000100110100_1000001001010101000;
        7'd26 : d = 31'b000101000000_1000001010000011100;
        7'd27 : d = 31'b000101001011_1000001010110011101;
        7'd28 : d = 31'b000101010111_1000001011100101010;
        7'd29 : d = 31'b000101100010_1000001100011000011;
        7'd30 : d = 31'b000101101110_1000001101001101001;
        7'd31 : d = 31'b000101111001_1000001110000011010;
        7'd32 : d = 31'b000110000100_1000001110111010111;
        7'd33 : d = 31'b000110010000_1000001111110100000;
        7'd34 : d = 31'b000110011011_1000010000101110100;
        7'd35 : d = 31'b000110100110_1000010001101010011;
        7'd36 : d = 31'b000110110001_1000010010100111101;
        7'd37 : d = 31'b000110111100_1000010011100110010;
        7'd38 : d = 31'b000111000111_1000010100100110001;
        7'd39 : d = 31'b000111010010_1000010101100111011;
        7'd40 : d = 31'b000111011101_1000010110101001110;
        7'd41 : d = 31'b000111101000_1000010111101101011;
        7'd42 : d = 31'b000111110010_1000011000110010001;
        7'd43 : d = 31'b000111111101_1000011001111000001;
        7'd44 : d = 31'b001000000111_1000011010111111001;
        7'd45 : d = 31'b001000010010_1000011100000111010;
        7'd46 : d = 31'b001000011100_1000011101010000011;
        7'd47 : d = 31'b001000100110_1000011110011010101;
        7'd48 : d = 31'b001000110001_1000011111100101110;
        7'd49 : d = 31'b001000111011_1000100000110001110;
        7'd50 : d = 31'b001001000101_1000100001111110110;
        7'd51 : d = 31'b001001001111_1000100011001100100;
        7'd52 : d = 31'b001001011001_1000100100011011001;
        7'd53 : d = 31'b001001100010_1000100101101010100;
        7'd54 : d = 31'b001001101100_1000100110111010101;
        7'd55 : d = 31'b001001110110_1000101000001011100;
        7'd56 : d = 31'b001001111111_1000101001011101000;
        7'd57 : d = 31'b001010001001_1000101010101111001;
        7'd58 : d = 31'b001010010010_1000101100000001110;
        7'd59 : d = 31'b001010011011_1000101101010101000;
        7'd60 : d = 31'b001010100100_1000101110101000101;
        7'd61 : d = 31'b001010101101_1000101111111100110;
        7'd62 : d = 31'b001010110110_1000110001010001011;
        7'd63 : d = 31'b001010111111_1000110010100110010;
        7'd64 : d = 31'b001011000111_1000110011111011011;
        7'd65 : d = 31'b001011010000_1000110101010000111;
        7'd66 : d = 31'b001011011000_1000110110100110100;
        7'd67 : d = 31'b001011100001_1000110111111100011;
        7'd68 : d = 31'b001011101001_1000111001010010010;
        7'd69 : d = 31'b001011110001_1000111010101000011;
        7'd70 : d = 31'b001011111001_1000111011111110011;
        7'd71 : d = 31'b001100000001_1000111101010100100;
        7'd72 : d = 31'b001100001001_1000111110101010100;
        7'd73 : d = 31'b001100010001_1001000000000000011;
        7'd74 : d = 31'b001100011000_1001000001010110000;
        7'd75 : d = 31'b001100100000_1001000010101011100;
        7'd76 : d = 31'b001100100111_1001000100000000110;
        7'd77 : d = 31'b001100101110_1001000101010101101;
        7'd78 : d = 31'b001100110101_1001000110101010001;
        7'd79 : d = 31'b001100111100_1001000111111110011;
        7'd80 : d = 31'b001101000011_1001001001010010000;
        7'd81 : d = 31'b001101001010_1001001010100101001;
        7'd82 : d = 31'b001101010000_1001001011110111110;
        7'd83 : d = 31'b001101010111_1001001101001001101;
        7'd84 : d = 31'b001101011101_1001001110011011000;
        7'd85 : d = 31'b001101100011_1001001111101011100;
        7'd86 : d = 31'b001101101001_1001010000111011011;
        7'd87 : d = 31'b001101101111_1001010010001010010;
        7'd88 : d = 31'b001101110101_1001010011011000011;
        7'd89 : d = 31'b001101111010_1001010100100101100;
        7'd90 : d = 31'b001110000000_1001010101110001110;
        7'd91 : d = 31'b001110000101_1001010110111100111;
        7'd92 : d = 31'b001110001011_1001011000000110111;
        7'd93 : d = 31'b001110010000_1001011001001111110;
        7'd94 : d = 31'b001110010101_1001011010010111100;
        7'd95 : d = 31'b001110011010_1001011011011110000;
        7'd96 : d = 31'b001110011110_1001011100100011001;
        7'd97 : d = 31'b001110100011_1001011101100110111;
        7'd98 : d = 31'b001110100111_1001011110101001011;
        7'd99 : d = 31'b001110101011_1001011111101010010;
        7'd100 : d = 31'b001110110000_1001100000101001101;
        7'd101 : d = 31'b001110110100_1001100001100111100;
        7'd102 : d = 31'b001110110111_1001100010100011110;
        7'd103 : d = 31'b001110111011_1001100011011110010;
        7'd104 : d = 31'b001110111111_1001100100010111001;
        7'd105 : d = 31'b001111000010_1001100101001110001;
        7'd106 : d = 31'b001111000101_1001100110000011011;
        7'd107 : d = 31'b001111001001_1001100110110110110;
        7'd108 : d = 31'b001111001100_1001100111101000001;
        7'd109 : d = 31'b001111001110_1001101000010111100;
        7'd110 : d = 31'b001111010001_1001101001000100111;
        7'd111 : d = 31'b001111010100_1001101001110000001;
        7'd112 : d = 31'b001111010110_1001101010011001010;
        7'd113 : d = 31'b001111011000_1001101011000000010;
        7'd114 : d = 31'b001111011010_1001101011100100111;
        7'd115 : d = 31'b001111011100_1001101100000111011;
        7'd116 : d = 31'b001111011110_1001101100100111011;
        7'd117 : d = 31'b001111100000_1001101101000101000;
        7'd118 : d = 31'b001111100001_1001101101100000001;
        7'd119 : d = 31'b001111100011_1001101101111000111;
        7'd120 : d = 31'b001111100100_1001101110001111000;
        7'd121 : d = 31'b001111100101_1001101110100010100;
        7'd122 : d = 31'b001111100110_1001101110110011100;
        7'd123 : d = 31'b001111100110_1001101111000001101;
        7'd124 : d = 31'b001111100111_1001101111001101001;
        7'd125 : d = 31'b000000000000_1001101111010101110;
        7'd126 : d = 31'b000000000000_1001101111011011101;
        7'd127 : d = 31'b000000000000_1001101111011110100;
        default: d = 31'd0;
        endcase
    end
    
    // Output Data
    always @(posedge clock) begin
        c1 <= d[30:19];
        c0 <= d[18:0];
    end    
endmodule
